// this file is immediate number generator for single cycle processor.
// ISA based on RV32I

module immgen (
    input [31:0] instruction,
    output reg [31:0] imm
);
    
endmodule